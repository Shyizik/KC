library verilog;
use verilog.vl_types.all;
entity function_f4_Yukhymchuk is
    port(
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        fnor_nor        : out    vl_logic;
        fnand_nand      : out    vl_logic
    );
end function_f4_Yukhymchuk;
