library verilog;
use verilog.vl_types.all;
entity testbench_demux_Yukhymchuk is
end testbench_demux_Yukhymchuk;
